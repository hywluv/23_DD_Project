`timescale 1ns / 1ps

module clk_vga( 
	input clk, 
	output reg clk_vga
);
	 
	reg [2:0] cnt;

	initial begin
		cnt = 32'b0;
	end

	wire[2:0] cnt_next;
	assign cnt_next = cnt + 1'b1;

	always @(posedge clk) begin
		if(cnt < 2)begin
			cnt <= cnt_next;
		end
		else begin
			cnt <= 0;
			clk_1s <= ~clk_1s;
		end
	end

endmodule
